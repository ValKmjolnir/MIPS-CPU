module hazard();



endmodule